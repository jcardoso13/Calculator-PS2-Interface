//
// VERSAT PROGRAM MEMORY DEFINES
//

// PROG address width
`define PROG_ADDR_W 9

// ROM address width
`define PROG_ROM_ADDR_W 4

// Program memory address width
`define PROG_RAM_ADDR_W 8

// Memory map
`define PROG_ROM `PROG_ADDR_W'h0
`define PROG_RAM `PROG_ADDR_W'h100

